library verilog;
use verilog.vl_types.all;
entity MiniMIPS_testbench is
end MiniMIPS_testbench;
