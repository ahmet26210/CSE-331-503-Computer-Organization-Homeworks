module mult32();








endmodule



